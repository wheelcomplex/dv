// <insert copyright notice here>

module main
